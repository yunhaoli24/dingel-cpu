LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX3 IS
PORT(
	I,BACK:IN STD_LOGIC;
	DATA,BIN,RIN:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	MUX3_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END MUX3;

ARCHITECTURE A OF MUX3 IS
BEGIN
    PROCESS
     BEGIN 
       IF(I='0') THEN     			
            MUX3_OUT<=DATA;
	   ELSIF(BACK='0')THEN 
			MUX3_OUT<=BIN;			
	   ELSE
			MUX3_OUT<=RIN;
		END IF;
    END PROCESS;
END A;


