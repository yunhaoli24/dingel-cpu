LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CONTROM IS
PORT(ADDR: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
     UA:OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
     O:OUT STD_LOGIC_VECTOR(20 DOWNTO 0)
    );
END CONTROM;
ARCHITECTURE A OF CONTROM IS
SIGNAL DATAOUT: STD_LOGIC_VECTOR(26 DOWNTO 0);
BEGIN 
    PROCESS
    BEGIN
        CASE ADDR IS    
        --        ΢��ַ                         ΢ָ��
            WHEN "000000" => DATAOUT<="110100100011111101100000000";--ȡ��ַ
            WHEN "000001" => DATAOUT<="100010100011111110000000000";--MOV
            WHEN "000010" => DATAOUT<="100010100010111011000000000";--IN
            WHEN "000011" => DATAOUT<="100011101101111111000000000";--DEC
            WHEN "000100" => DATAOUT<="100001100111111111000000000";--TEST
            WHEN "000101" => DATAOUT<="100000100011111111010000000";--JB
            WHEN "000110" => DATAOUT<="100000100011111111001000000";--JZ
            WHEN "000111" => DATAOUT<="010000100011111110000000000";--JMP
            WHEN "001000" => DATAOUT<="100001100111111111000000000";--CMP
            WHEN "001001" => DATAOUT<="100011100001111111000000000";--ADD
            WHEN "001010" => DATAOUT<="100000000011011111000000000";--OUT
            WHEN "001011" => DATAOUT<="101000000011111111000001100";--LAD
            WHEN "001100" => DATAOUT<="100010100011111011000000000";--LAD2
            WHEN "001101" => DATAOUT<="101000111101111111000001110";--STO
            WHEN "001110" => DATAOUT<="100000000011101111000000000";--STO2
            WHEN "001111" => DATAOUT<="100011101001111111000000000";--INC

            WHEN "100000" => DATAOUT<="010000100011111110000000000";--jb
            WHEN "010000" => DATAOUT<="010000100011111110000000000";--jz

            WHEN OTHERS   => DATAOUT<="110100100011111101100000000";
        END CASE;
        UA(5 DOWNTO 0)<=DATAOUT(5 DOWNTO 0);
        O(20 DOWNTO 0)<=DATAOUT(26 DOWNTO 6);
    END PROCESS;
END A;


