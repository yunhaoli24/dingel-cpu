LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PSW IS
PORT(
     C,Z,LDPSW: IN STD_LOGIC;
     CF,ZF: OUT STD_LOGIC
    );
END PSW;

ARCHITECTURE A OF PSW IS
BEGIN 
     PROCESS(LDPSW)
     BEGIN
         IF(LDPSW'EVENT AND LDPSW='1') THEN
             CF<=C;
             ZF<=Z;
         END IF;
     END PROCESS;
END A;


