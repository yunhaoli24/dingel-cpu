LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY F3 IS 
PORT(
    D:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    UA3,UA2,UA1,UA0: OUT STD_LOGIC
    );
END F3;
ARCHITECTURE A OF F3 IS
BEGIN
    UA3<=D(3);
    UA2<=D(2);
    UA1<=D(1);
    UA0<=D(0);
END A;




