LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MODE_CONTROL IS
PORT(
	CF,ZF:IN STD_LOGIC;
	T1,T2,T3,T4,CLR:IN STD_LOGIC;
	DIN:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLK:IN STD_LOGIC;
	LOAD,LDPC,LDAR,LDIR,LDRI,RD_B,RS_B,S1,S0:OUT STD_LOGIC;
	ALU_B,LDAC,LDDR,CS_I,SW_B,LED_B,LDPSW:OUT STD_LOGIC
	);
END MODE_CONTROL;
ARCHITECTURE A OF MODE_CONTROL IS
SIGNAL YIMA:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL IN1,MOV,CMP,JB,ADD,INC,JMP,OUT1:STD_LOGIC;
SIGNAL M:STD_LOGIC:='0';
BEGIN
	P1:PROCESS(CLR,T4)
	BEGIN
		IF(CLR='0')THEN
			M<='0';
		ELSIF(T4'EVENT AND T4='0')THEN
			M<=NOT M;
		END IF;
	END PROCESS P1;
	P2:PROCESS(CLK)
	BEGIN
		CASE DIN(3 DOWNTO 0)IS
			WHEN "0000"=>YIMA<="00000001";
			WHEN "0001"=>YIMA<="00000010";
			WHEN "0010"=>YIMA<="00000100";
			WHEN "0011"=>YIMA<="00001000";
			WHEN "0100"=>YIMA<="00010000";
			WHEN "0101"=>YIMA<="00100000";
			WHEN "0110"=>YIMA<="01000000";
			WHEN "0111"=>YIMA<="10000000";
			WHEN OTHERS=>YIMA<="00000000";
		END CASE;
		LOAD<=NOT((JMP AND T4 AND (NOT M)) OR (JB AND T4 AND (NOT M) AND (CF AND (NOT ZF))));
		
		LDPC<=(T1 AND (NOT CLK) AND (NOT M)) 
				OR (( MOV OR JB OR JMP) AND T3 AND (NOT CLK) AND (NOT M)) 
				OR (JB AND T4 AND (NOT CLK) AND (NOT M) AND (CF AND (NOT ZF))) 
				OR (JMP AND T4 AND (NOT CLK) AND (NOT M));
				
		LDAR<=(T1 OR ((MOV OR JB OR JMP) AND T3)) AND (NOT CLK) AND (NOT M);

		LDIR<=T2 AND (NOT CLK) AND (NOT M);
		
		LDRI<=(IN1 AND T3 AND (NOT CLK) AND (NOT M))
				OR (MOV AND T4 AND (NOT CLK) AND (NOT M))
				OR (ADD AND T1 AND (NOT CLK) AND M)
				OR (INC AND T4 AND (NOT CLK) AND (NOT M));

		RD_B<=NOT(
					(CMP AND T4 AND (NOT M))
					OR (ADD AND T4 AND (NOT M))
					OR (INC AND T3 AND (NOT M))
				);

		RS_B<=NOT((CMP OR ADD OR OUT1) AND T3 AND (NOT M));

		S1<=INC AND T4 AND (NOT M);

		S0<=CMP AND T1 AND M;

		ALU_B<=NOT((ADD AND T1 AND M) OR (INC AND T4 AND (NOT M)));
		
		LDAC<=(CMP OR ADD OR INC) AND T3 AND (NOT CLK) AND (NOT M);
		
		LDDR<=(CMP OR ADD) AND T4 AND (NOT CLK) AND (NOT M);
		
		CS_I<=NOT(
				(T2 AND (NOT M) OR (MOV AND T4 AND (NOT M))
				OR (JB AND T4 AND (NOT M) AND (CF AND (NOT ZF)))
				OR (JMP AND T4 AND (NOT M))
				);

		SW_B<=NOT(IN1 AND T3 AND (NOT M));

		LED_B<=NOT(IN1 AND T3 AND (NOT M));

		LDPSW<=CMP AND T1 AND (NOT CLK) AND M;
	END PROCESS P2;
	OUT1<=YIMA(7);
	JMP<=YIMA(6);
	INC<=YIMA(5);
	ADD<=YIMA(4);
	JB<=YIMA(3);
	CMP<=YIMA(2);
	MOV<=YIMA(1);
	IN1<=YIMA(0);
END A;
