LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ROM IS 
PORT(
	DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDR:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	CS_I:IN STD_LOGIC
);
END ROM;
ARCHITECTURE A OF ROM IS

--  ע�Ƿ���    ָ���ʽ(OP)    Rs Rd     addr   
--    MOV            0001       XX Rd    XXXXXXXX
--    INT            0010       XX Rd    XXXXXXXX
--    TEST           0011       Rs XX    XXXXXXXX
--    JB             0100       XX XX     addr
--    MUL            0101       Rs Rd    XXXXXXXX
--    ADD            0110       Rs Rd    XXXXXXXX
--    DEC            0111       XX Rd    XXXXXXXX
--    JZ             1000       XX XX     addr
--    OUT            1001       Rs XX    XXXXXXXX
--    JMP            1010       XX XX     addr
BEGIN
	DOUT<="0001000100000010" WHEN ADDR="00000000" AND CS_I='0' ELSE--MOV R1,2H
          "0001001000000110" WHEN ADDR="00000001" AND CS_I='0' ELSE--MOV R2,6H
          "0001001100000111" WHEN ADDR="00000010" AND CS_I='0' ELSE--MOV R3,7H
          "0001000000000011" WHEN ADDR="00000011" AND CS_I='0' ELSE--MOV R0,3H

		  "0000000000000000";
END A;


