LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ROM IS
PORT(
		DOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		ADDR:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		CS:IN STD_LOGIC
);
END ROM;
ARCHITECTURE A OF ROM IS
BEGIN
	DOUT<=	"10000000" WHEN ADDR="00000000" AND CS='0' ELSE
			"10010001" WHEN ADDR="00000001" AND CS='0' ELSE
			"00000001" WHEN ADDR="00000010" AND CS='0' ELSE
			"10010010" WHEN ADDR="00000011" AND CS='0' ELSE
			"00000000" WHEN ADDR="00000100" AND CS='0' ELSE
			"10100001" WHEN ADDR="00000101" AND CS='0' ELSE
			"10110000" WHEN ADDR="00000110" AND CS='0' ELSE
			"00001101" WHEN ADDR="00000111" AND CS='0' ELSE
			"11000110" WHEN ADDR="00001000" AND CS='0' ELSE
			"11010001" WHEN ADDR="00001001" AND CS='0' ELSE
			"11010001" WHEN ADDR="00001010" AND CS='0' ELSE
			"11100000" WHEN ADDR="00001011" AND CS='0' ELSE
			"10000101" WHEN ADDR="00001100" AND CS='0' ELSE
			"11111000" WHEN ADDR="00001101" AND CS='0' ELSE
			"11100000" WHEN ADDR="00001110" AND CS='0' ELSE
			"00001101" WHEN ADDR="00001111" AND CS='0' ELSE
			"00000000";
END A;


