LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONVERT IS
PORT(
	IRCODE:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	OP:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	I3,I2,I1,I0:OUT STD_LOGIC
);
END CONVERT;
ARCHITECTURE A OF CONVERT IS
BEGIN
	OP<=IRCODE(7 DOWNTO 4);
	I3<=IRCODE(3);
	I2<=IRCODE(2);
	I1<=IRCODE(1);
	I0<=IRCODE(0);
END A;
