LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ROM IS 
PORT(
	DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDR:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	CS_I:IN STD_LOGIC
);
END ROM;
ARCHITECTURE A OF ROM IS

--  ע�Ƿ���    ָ���ʽ(OP)    Rs Rd     addr
   
--    MOV           0001        XX Rd     im

--    IN            0010        XX Rd    XXXXXXXX

--    DEC           0011        XX Rd    XXXXXXXX

--    TEST          0100        XX Rd     addr

--    JB            0101        XX XX     addr

--    JZ            0110        XX XX     addr

--    JMP           0111        XX XX     addr

--    CMP           1000        Rs Rd    XXXXXXXX

--    ADD           1001        Rs Rd    XXXXXXXX

--    OUT           1010        Rs XX    XXXXXXXX

--    LAD           1011        Rs(Rd)   XXXXXXXX

--    STO           1101        Rs(Rd)   XXXXXXXX

--    INC           1111        XX Rd    XXXXXXXX

BEGIN
	--DOUT<="0001000000000000" WHEN ADDR="00000000" AND CS_I='0' ELSE--MOV R0,0H
          --"0001000100000101" WHEN ADDR="00000001" AND CS_I='0' ELSE--MOV R1,5H
          --"0010001000000000" WHEN ADDR="00000010" AND CS_I='0' ELSE--FLAG1:IN R2
          --"1101100000000000" WHEN ADDR="00000011" AND CS_I='0' ELSE--STO R2,(R0)
          --"1111000000000000" WHEN ADDR="00000100" AND CS_I='0' ELSE--INC R0
          --"1000000100000000" WHEN ADDR="00000101" AND CS_I='0' ELSE--CMP R0,R1
          --"0110000000001000" WHEN ADDR="00000110" AND CS_I='0' ELSE--JZ FLAG2
          --"0111000000000010" WHEN ADDR="00000111" AND CS_I='0' ELSE--JMP FLAG1
          --"0001001100000101" WHEN ADDR="00001000" AND CS_I='0' ELSE--FLAG2:MOV R3,05H
          --"1101110000000000" WHEN ADDR="00001001" AND CS_I='0' ELSE--STO R3,(R0)
															---------����10����
	DOUT<="0001000000000000" WHEN ADDR="00000000" AND CS_I='0' ELSE--MOV R0,0H
          "0001000100001010" WHEN ADDR="00000001" AND CS_I='0' ELSE--MOV R1,10
          "0010001000000000" WHEN ADDR="00000010" AND CS_I='0' ELSE--FLAG1:IN R2
          "1101100000000000" WHEN ADDR="00000011" AND CS_I='0' ELSE--STO R2,(R0)
          "1111000000000000" WHEN ADDR="00000100" AND CS_I='0' ELSE--INC R0
          "1000000100000000" WHEN ADDR="00000101" AND CS_I='0' ELSE--CMP R0,R1
          "0101000000000010" WHEN ADDR="00000110" AND CS_I='0' ELSE--JB FLAG1
															---------��ʼ������
          "0001000100010100" WHEN ADDR="00000111" AND CS_I='0' ELSE--MOV R1,20
          "0001001000000001" WHEN ADDR="00001000" AND CS_I='0' ELSE--MOV R2,1H
          "1101100000000000" WHEN ADDR="00001001" AND CS_I='0' ELSE--FLAG2:ST0 R2,(R0)
          "1111000000000000" WHEN ADDR="00001010" AND CS_I='0' ELSE--INC R0
          "1000000100000000" WHEN ADDR="00001011" AND CS_I='0' ELSE--CMP R0,R1
          "0101000000001001" WHEN ADDR="00001100" AND CS_I='0' ELSE--JB FALG2
															---------��¼����
          "0001000100000000" WHEN ADDR="00001101" AND CS_I='0' ELSE--MOV R1,0H
          "0001000000000001" WHEN ADDR="00001110" AND CS_I='0' ELSE--FLAG3:MOV R0,1H
          "1001010000000000" WHEN ADDR="00001111" AND CS_I='0' ELSE--ADD RO,R1
          "1011011000000000" WHEN ADDR="00010000" AND CS_I='0' ELSE--FLAG4:LAD (R1),R2
          "1011001100000000" WHEN ADDR="00010001" AND CS_I='0' ELSE--LAD (R0),R3
          "1000101100000000" WHEN ADDR="00010010" AND CS_I='0' ELSE--CMP R2,R3
          "0110000000011100" WHEN ADDR="00010011" AND CS_I='0' ELSE--JZ ADD_ONE
          "1111000000000000" WHEN ADDR="00010100" AND CS_I='0' ELSE--FLAG5:INC RO
          "0001001000001010" WHEN ADDR="00010101" AND CS_I='0' ELSE--MOV R2,10
          "1000001000000000" WHEN ADDR="00010110" AND CS_I='0' ELSE--CMP R0,R2
          "0101000000010000" WHEN ADDR="00010111" AND CS_I='0' ELSE--JB FLAG4
          "1111000100000000" WHEN ADDR="00011000" AND CS_I='0' ELSE--INC R1
          "1000011000000000" WHEN ADDR="00011001" AND CS_I='0' ELSE--CMP R1,R2
          "0101000100001110" WHEN ADDR="00011010" AND CS_I='0' ELSE--JB FLAG3
          "0111000000100110" WHEN ADDR="00011011" AND CS_I='0' ELSE--JMP FALG6
          "0001001100011111" WHEN ADDR="00011100" AND CS_I='0' ELSE--ADD_ONE:MOV R3,31
          "1101011100000000" WHEN ADDR="00011101" AND CS_I='0' ELSE--STO R1,(R3)
          "0001001100001010" WHEN ADDR="00011110" AND CS_I='0' ELSE--MOV R3,10

          "1001110100000000" WHEN ADDR="00011111" AND CS_I='0' ELSE--ADD R1,R3
          "1011011100000000" WHEN ADDR="00100000" AND CS_I='0' ELSE--LAD (R1),R3
          "1111001100000000" WHEN ADDR="00100001" AND CS_I='0' ELSE--INC R3
          "1101110100000000" WHEN ADDR="00100010" AND CS_I='0' ELSE--STO R3,(R1)
          "0001001100011111" WHEN ADDR="00100011" AND CS_I='0' ELSE--MOV R3,31
          "1011110100000000" WHEN ADDR="00100100" AND CS_I='0' ELSE--LAD (R3),R1
          "0111000000010100" WHEN ADDR="00100101" AND CS_I='0' ELSE--JMP FALG5

          "0001000000000000" WHEN ADDR="00100110" AND CS_I='0' ELSE--FALG6:MOV R0,0
          "0001000100010100" WHEN ADDR="00100111" AND CS_I='0' ELSE--MOV R1,20
          "0001001000011101" WHEN ADDR="00101000" AND CS_I='0' ELSE--MOV R2,29
          "1011001100000000" WHEN ADDR="00101001" AND CS_I='0' ELSE--LAD (R0),R3
          "1101111000000000" WHEN ADDR="00101010" AND CS_I='0' ELSE--STO R3,(R2)
          "1111001000000000" WHEN ADDR="00101011" AND CS_I='0' ELSE--INC R2
          "0001001100001010" WHEN ADDR="00101100" AND CS_I='0' ELSE--MOV R3,10
          "1001110000000000" WHEN ADDR="00101101" AND CS_I='0' ELSE--ADD R0,R3
          "1011001100000000" WHEN ADDR="00101110" AND CS_I='0' ELSE--LAD (R0),R3
          "1101111000000000" WHEN ADDR="00101111" AND CS_I='0' ELSE--STO R3,(R2)
          "0001000000000000" WHEN ADDR="00110000" AND CS_I='0' ELSE--MOV R0,0
          "1111000000000000" WHEN ADDR="00110001" AND CS_I='0' ELSE--FLAG7:INC R0
          "0001000100001010" WHEN ADDR="00110010" AND CS_I='0' ELSE--MOV R1,10
          "1001000100000000" WHEN ADDR="00110011" AND CS_I='0' ELSE--ADD R1,R0
          "1011011000000000" WHEN ADDR="00110100" AND CS_I='0' ELSE--LAD (R1),R2
          "1000111000000000" WHEN ADDR="00110101" AND CS_I='0' ELSE--CMP R3,R2
          "0101000000111011" WHEN ADDR="00110110" AND CS_I='0' ELSE--JB SAVE

          "0001000100001001" WHEN ADDR="00110111" AND CS_I='0' ELSE--MOV R1,9
          "1000000100000000" WHEN ADDR="00111000" AND CS_I='0' ELSE--CMP R0,R1
          "0101000000110001" WHEN ADDR="00111001" AND CS_I='0' ELSE--JB FLAG7
          "0111000001000100" WHEN ADDR="00111010" AND CS_I='0' ELSE--JMP END

          "0001000100011110" WHEN ADDR="00111011" AND CS_I='0' ELSE--SAVE:MOV R1,30
          "1101100100000000" WHEN ADDR="00111100" AND CS_I='0' ELSE--STO R2,(R1)
          "1011011100000000" WHEN ADDR="00111101" AND CS_I='0' ELSE--LAD (R1),R3
          "1011001000000000" WHEN ADDR="00111110" AND CS_I='0' ELSE--LAD (R0),R2
          "0001000100011101" WHEN ADDR="00111111" AND CS_I='0' ELSE--MOV R1,29
          "1101100100000000" WHEN ADDR="01000000" AND CS_I='0' ELSE--STO R2,(R1)
          "0001000100001001" WHEN ADDR="01000001" AND CS_I='0' ELSE--MOV R1,9
          "1000000100000000" WHEN ADDR="01000010" AND CS_I='0' ELSE--CMP R0,R1
          "0101000000110001" WHEN ADDR="01000011" AND CS_I='0' ELSE--JB FLAG7

          "0001000000011101" WHEN ADDR="01000100" AND CS_I='0' ELSE--END:MOV R0,29
          "1011100000000000" WHEN ADDR="01000101" AND CS_I='0' ELSE--LAD R2,(R0)
          "1111000000000000" WHEN ADDR="01000110" AND CS_I='0' ELSE--INC R0
          "1011110000000000" WHEN ADDR="01000111" AND CS_I='0' ELSE--LAD R3,(R0)
          "1010100000000000" WHEN ADDR="01001000" AND CS_I='0' ELSE--OUT R2
          "1010110000000000" WHEN ADDR="01001001" AND CS_I='0' ELSE--OUT R3
          --"1011011000000000" WHEN ADDR="00010000" AND CS_I='0' ELSE--FLAG4:LAD (R1),R2
          --"1111000000000000" WHEN ADDR="00010001" AND CS_I='0' ELSE--INC R0
          --"0001001100011111" WHEN ADDR="00010010" AND CS_I='0' ELSE--MOV R3,31
          --"1101001100000000" WHEN ADDR="00010011" AND CS_I='0' ELSE--STO R0,(R3)
          --"1011001100000000" WHEN ADDR="00010100" AND CS_I='0' ELSE--LAD (R0),R3
          --"1000101100000000" WHEN ADDR="00010101" AND CS_I='0' ELSE--CMP R2,R3

          --"0110000000011110" WHEN ADDR="00010110" AND CS_I='0' ELSE--JZ FLAG6
          --"0001001100001001" WHEN ADDR="00010111" AND CS_I='0' ELSE--MOV R3,09H
          --"1000001100000000" WHEN ADDR="00011000" AND CS_I='0' ELSE--CMP R0,R3
          --"0101000000010000" WHEN ADDR="00011001" AND CS_I='0' ELSE--JB FLAG4

          --"1111000100000000" WHEN ADDR="00011010" AND CS_I='0' ELSE--FLAG5:INC R1
          --"1111001100000000" WHEN ADDR="00011011" AND CS_I='0' ELSE--INC R3
          --"1000011100000000" WHEN ADDR="00011100" AND CS_I='0' ELSE--CMP R1,R3
          --"0101000000001110" WHEN ADDR="00011101" AND CS_I='0' ELSE--JB FLAG3
          --"0111000000101011" WHEN ADDR="00011110" AND CS_I='0' ELSE--JMP FLAG7
          --"0001001000001010" WHEN ADDR="00011111" AND CS_I='0' ELSE--FLAG6:MOV R2,10H
          --"0001000000000000" WHEN ADDR="00100000" AND CS_I='0' ELSE--MOV R0,0H
          --"1001010000000000" WHEN ADDR="00100001" AND CS_I='0' ELSE--ADD R0,R1
          --"1001100000000000" WHEN ADDR="00100010" AND CS_I='0' ELSE--ADD R0,R2
          --"1011001100000000" WHEN ADDR="00100011" AND CS_I='0' ELSE--LAD (R0),R3
          --"1111001100000000" WHEN ADDR="00100100" AND CS_I='0' ELSE--INC R3
          --"1101110000000000" WHEN ADDR="00100101" AND CS_I='0' ELSE--STO R3,(R0)
          --"0001001100011111" WHEN ADDR="00100110" AND CS_I='0' ELSE--MOV R3,31
          --"1011110000000000" WHEN ADDR="00100111" AND CS_I='0' ELSE--LAD (R3),R0

          --"0001001100001001" WHEN ADDR="00101000" AND CS_I='0' ELSE--MOV R3,09H
          --"1000001100000000" WHEN ADDR="00101001" AND CS_I='0' ELSE--CMP R0,R3
          --"0101000000010000" WHEN ADDR="00101010" AND CS_I='0' ELSE--JB FLAG4

          --"0111000000011010" WHEN ADDR="00101011" AND CS_I='0' ELSE--JMP FLAG5
          --"0001000100000001" WHEN ADDR="00101100" AND CS_I='0' ELSE--FLAG7:MOV R1,1H
          --"0001001000000100" WHEN ADDR="00101101" AND CS_I='0' ELSE--MOV R2,4H
          --"1010010000000000" WHEN ADDR="00101110" AND CS_I='0' ELSE--OUT R1
          --"1010100000000000" WHEN ADDR="00101111" AND CS_I='0' ELSE--OUT R2
          --"1111000000000000" WHEN ADDR="00000101" AND CS_I='0' ELSE--
          --"1000000100000000" WHEN ADDR="00000110" AND CS_I='0' ELSE--
          --"0101000000000100" WHEN ADDR="00000111" AND CS_I='0' ELSE--
          --"1010110000000000" WHEN ADDR="00001000" AND CS_I='0' ELSE--
          --"0001000000000011" WHEN ADDR="00000110" AND CS_I='0' ELSE--
          --"0001001000000110" WHEN ADDR="00000100" AND CS_I='0' ELSE--
          --"0001001100000111" WHEN ADDR="00000101" AND CS_I='0' ELSE--
		  "0000000000000000";
END A;
