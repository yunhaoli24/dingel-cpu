LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ADDR IS 
PORT(
     I15,I14,I13,I12:IN STD_LOGIC;
     ZF,CF,T4,P1,P2:IN STD_LOGIC;
     SE5,SE4,SE3,SE2,SE1,SE0:OUT STD_LOGIC
);
END ADDR;
ARCHITECTURE A OF ADDR IS
BEGIN
     SE5<=NOT( NOT(CF) AND P2 AND T4);
     SE4<='1'; 
     SE3<=NOT(I15 AND P1 AND T4);
     SE2<=NOT(I14 AND P1 AND T4);
     SE1<=NOT(I13 AND P1 AND T4);
     SE0<=NOT(I12 AND P1 AND T4);
END A;


